
module serial_crc_ccitt (
sys_clk     ,
sys_resetb   ,
enable  ,
//init    , 
data_in ,
CMD, 
CRC_M,
init,

CTS,
CTS_error
);
//-----------Input Ports---------------
input        sys_clk;
input        sys_resetb;
input        enable;              // ?��?��?�� -> shift마다 발생 
//input init    ;
input       data_in;             // 1비트?�� ?��?��
input [3:0] CMD;
input [3:0] CRC_M;         // ?��?��?�� ?��맷의 CRC ?��?���?
input       init;          // ?��?��?�� ?��맷이 종료?��?�� ?��?��?��?�� 1
//-----------Output Ports---------------
output       CTS;          // Clear To Send
output       CTS_error;    // Clear To Send ?���? CRC값이 맞�? ?��?��
//------------Internal Variables--------
reg  [3:0] lfsr;
reg  [2:0] count_init;
reg        flag;
reg  [3:0] enable_counter;
reg        report_flag;
reg  [5:0] count_enable;

wire [3:0] crc_out;
//-------------Code Start-----------------
assign crc_out = lfsr;
assign CTS           = (init==1'b1&&crc_out==CRC_M)? 1'b1 : 1'b0; // ?��?��?�� ?��맷이 종료?��?�� ?��?��?��?�� Clear To Send
assign CTS_error     = (init==1'b1&&crc_out!=CRC_M)? 1'b1 : 1'b0; // ?��?��?�� ?��맷이 종료?��?�� ?��?��?��?�� Clear To Send Error(CRC�? 불일�?)
// Logic to CRC Calculation
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
always @ (posedge sys_clk or negedge sys_resetb)
if (!sys_resetb) begin
  lfsr <= 4'b0000;
end 
else if (init) begin
  lfsr <= 4'b0000;
end
else if (enable==1'b1&&flag==1'b1&&!report_flag&&enable_counter<4'h8) begin // enable == shift, CRC_M �?분�? ?��?��?���? ?��?��?�� ?��(flag==1'b1),enable_counter -> 1 byte(0~7) calculate
    lfsr[0]  <= data_in ^ lfsr[3];                            // ?��?���? 같이 CRC-4-ITU�? ?��?��?��?���? 계산
    lfsr[1]  <= lfsr[0] ^ data_in ^ lfsr[3];
    lfsr[2]  <= lfsr[1];
    lfsr[3]  <= lfsr[2];
end 

always@(posedge sys_clk or negedge sys_resetb) begin
  if(!sys_resetb) begin
    report_flag <= 1'b0;
  end
  else if(count_enable==5'd17) begin
    report_flag <= 1'b0;
  end  
  else if(CMD==4'b1110&&init)begin
    report_flag <= 1'b1;
  end
end

always@(posedge sys_clk or negedge sys_resetb) begin
  if(!sys_resetb) begin
    count_enable <= 5'b0;
  end
  else if(report_flag==1'b1&&enable) begin
    count_enable <= count_enable + 1'b1;
  end  
  else if(count_enable==5'd17) begin
    count_enable <= 5'b0;
  end
  else begin
    count_enable <= count_enable;
  end
end

////////////////////////////////////////////////////////////////////////////////////////////////
always @ (posedge sys_clk or negedge sys_resetb)begin
if (!sys_resetb) begin
  flag <= 1'b0;
  count_init <= 1'b1;
end
else if (init) begin
  flag <= 1'b0;
  count_init <= 3'd1;
end
else if(report_flag) begin
  count_init <= 3'b1;
end
else if (enable==1'b1&&flag==1'b0) begin
  count_init <= count_init + 1'b1;
  if(count_init==3'd4) begin
    flag <= 1'b1;
  end
end
end
////////////////////////////////////////////////////////////////////////////////////////////////{CRC_M,CMD} ?��?��?�� ?��맷의 첫번�? Byte?��?�� 4�? Bit�? 무시?���? ?��?�� 구현
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
always @ (posedge sys_clk or negedge sys_resetb)
begin
if (!sys_resetb) begin
    enable_counter <= 1'b0;
end
else if(init)
    enable_counter <= 1'b0;
else if(report_flag)
    enable_counter <= 4'b0;    
else if(enable) begin
    enable_counter <= enable_counter + 1'b1;
    if(enable_counter==4'd8)
       enable_counter <= 1'b0; 
end
else
    enable_counter <= enable_counter;
end
//8bit�? ?��?��, enable_counter -> 8?��?�� 0?���? 초기?��


///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
endmodule